//~~~~NEXT_PC_CALCULATION~~~//
`define PC_IF 2'b00
`define PC_EX 2'b01
`define PC_REG 2'b11
//~~~~~~~~~~~~~~~~~~~~~~~~~~//
