//~~~ALU CODES~~~//
`define ALU_ADD  4'b00_00
`define ALU_SUB  4'b00_01
`define ALU_AND  4'b01_00
`define ALU_OR   4'b01_01
`define ALU_XOR  4'b01_10
`define ALU_SHL  4'b10_00
`define ALU_SHR  4'b10_10
`define ALU_SHA  4'b10_11
`define ALU_SLT  4'b11_00
`define ALU_SLTU 4'b11_01
`define ALU_SRC1 4'b01_11
`define ALU_SRC2 4'b11_11
